library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package config is
	constant num_microsteps		:natural;
	type power_table_type is array (0 to 256) of natural range 0 to 1000;
	constant power_table		:power_table_type;
end package;

package body config is
	constant num_microsteps		:natural	:=	1;
	
	-- Power table: holds the values of a quarter sine wave, in 0.1%
	constant power_table		:power_table_type	:= (
		1000,	1000,	1000,	1000,	1000,	1000,	999,	999,
		999,	998,	998,	998,	997,	997,	996,	996,
		995,	995,	994,	993,	992,	992,	991,	990,
		989,	988,	987,	986,	985,	984,	983,	982,
		981,	980,	978,	977,	976,	974,	973,	972,
		970,	969,	967,	965,	964,	962,	960,	959,
		957,	955,	953,	951,	950,	948,	946,	944,
		942,	939,	937,	935,	933,	931,	929,	926,
		924,	922,	919,	917,	914,	912,	909,	907,
		904,	901,	899,	896,	893,	890,	888,	885,
		882,	879,	876,	873,	870,	867,	864,	861,
		858,	855,	851,	848,	845,	842,	838,	835,
		831,	828,	825,	821,	818,	814,	810,	807,
		803,	800,	796,	792,	788,	785,	781,	777,
		773,	769,	765,	761,	757,	753,	749,	741,
		745,	737,	733,	728,	724,	720,	716,	711,
		707,	703,	698,	694,	690,	685,	681,	676,
		672,	667,	662,	658,	653,	649,	644,	639,
		634,	630,	625,	620,	615,	610,	606,	601,
		596,	591,	586,	581,	576,	571,	566,	561,
		556,	550,	545,	540,	535,	530,	525,	519,
		514,	509,	504,	498,	493,	488,	482,	477,
		471,	466,	461,	455,	450,	444,	439,	433,
		428,	422,	416,	411,	405,	400,	394,	388,
		383,	377,	371,	366,	360,	354,	348,	343,
		337,	331,	325,	320,	314,	308,	302,	296,
		290,	284,	279,	273,	267,	261,	255,	249,
		243,	237,	231,	225,	219,	213,	207,	201,
		195,	189,	183,	177,	171,	165,	159,	153,
		147,	141,	135,	128,	122,	116,	110,	104,
		98,	92,	86,	80,	74,	67,	61,	55,
		49,	43,	37,	31,	25,	18,	12,	6,
		0
	);
end config;


