library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package config is
    constant num_microsteps     :natural;
   
end package;

package body config is
    constant num_microsteps     :natural    :=  1;
    

end config;


